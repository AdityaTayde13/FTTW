module thruwire(i_sw, o_led);
	input i_sw;
	output o_led;

	assign o_led = i_sw;
endmodule
